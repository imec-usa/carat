`timescale 1ns/1ps

// 32-bit Carry-Lookahead Adder (CLA)
// Flattened for synthesis - no hierarchical modules

module adder_32bit (
    input wire [31:0] a,
    input wire [31:0] b,
    output wire [31:0] sum
);

    // Propagate and Generate signals
    wire [31:0] p, g;

    // Carry signals
    wire [32:0] c;
    assign c[0] = 1'b0;

    // Block-level propagate and generate (8 blocks of 4 bits each)
    wire [7:0] block_p, block_g;
    wire [8:0] block_c;
    assign block_c[0] = 1'b0;

    // Generate P and G for all 32 bits
    assign p = a ^ b;  // Propagate
    assign g = a & b;  // Generate

    // =========================================================================
    // Block 0: bits [3:0]
    // =========================================================================
    // Carry chain
    assign c[1] = g[0] | (p[0] & c[0]);
    assign c[2] = g[1] | (p[1] & c[1]);
    assign c[3] = g[2] | (p[2] & c[2]);
    assign c[4] = g[3] | (p[3] & c[3]);

    // Block propagate and generate
    assign block_p[0] = p[0] & p[1] & p[2] & p[3];
    assign block_g[0] = g[3] | (p[3] & g[2]) | (p[3] & p[2] & g[1]) | (p[3] & p[2] & p[1] & g[0]);

    // =========================================================================
    // Block 1: bits [7:4]
    // =========================================================================
    assign c[5] = g[4] | (p[4] & c[4]);
    assign c[6] = g[5] | (p[5] & c[5]);
    assign c[7] = g[6] | (p[6] & c[6]);
    assign c[8] = g[7] | (p[7] & c[7]);

    assign block_p[1] = p[4] & p[5] & p[6] & p[7];
    assign block_g[1] = g[7] | (p[7] & g[6]) | (p[7] & p[6] & g[5]) | (p[7] & p[6] & p[5] & g[4]);

    // =========================================================================
    // Block 2: bits [11:8]
    // =========================================================================
    assign c[9]  = g[8]  | (p[8]  & c[8]);
    assign c[10] = g[9]  | (p[9]  & c[9]);
    assign c[11] = g[10] | (p[10] & c[10]);
    assign c[12] = g[11] | (p[11] & c[11]);

    assign block_p[2] = p[8] & p[9] & p[10] & p[11];
    assign block_g[2] = g[11] | (p[11] & g[10]) | (p[11] & p[10] & g[9]) | (p[11] & p[10] & p[9] & g[8]);

    // =========================================================================
    // Block 3: bits [15:12]
    // =========================================================================
    assign c[13] = g[12] | (p[12] & c[12]);
    assign c[14] = g[13] | (p[13] & c[13]);
    assign c[15] = g[14] | (p[14] & c[14]);
    assign c[16] = g[15] | (p[15] & c[15]);

    assign block_p[3] = p[12] & p[13] & p[14] & p[15];
    assign block_g[3] = g[15] | (p[15] & g[14]) | (p[15] & p[14] & g[13]) | (p[15] & p[14] & p[13] & g[12]);

    // =========================================================================
    // Block 4: bits [19:16]
    // =========================================================================
    assign c[17] = g[16] | (p[16] & c[16]);
    assign c[18] = g[17] | (p[17] & c[17]);
    assign c[19] = g[18] | (p[18] & c[18]);
    assign c[20] = g[19] | (p[19] & c[19]);

    assign block_p[4] = p[16] & p[17] & p[18] & p[19];
    assign block_g[4] = g[19] | (p[19] & g[18]) | (p[19] & p[18] & g[17]) | (p[19] & p[18] & p[17] & g[16]);

    // =========================================================================
    // Block 5: bits [23:20]
    // =========================================================================
    assign c[21] = g[20] | (p[20] & c[20]);
    assign c[22] = g[21] | (p[21] & c[21]);
    assign c[23] = g[22] | (p[22] & c[22]);
    assign c[24] = g[23] | (p[23] & c[23]);

    assign block_p[5] = p[20] & p[21] & p[22] & p[23];
    assign block_g[5] = g[23] | (p[23] & g[22]) | (p[23] & p[22] & g[21]) | (p[23] & p[22] & p[21] & g[20]);

    // =========================================================================
    // Block 6: bits [27:24]
    // =========================================================================
    assign c[25] = g[24] | (p[24] & c[24]);
    assign c[26] = g[25] | (p[25] & c[25]);
    assign c[27] = g[26] | (p[26] & c[26]);
    assign c[28] = g[27] | (p[27] & c[27]);

    assign block_p[6] = p[24] & p[25] & p[26] & p[27];
    assign block_g[6] = g[27] | (p[27] & g[26]) | (p[27] & p[26] & g[25]) | (p[27] & p[26] & p[25] & g[24]);

    // =========================================================================
    // Block 7: bits [31:28]
    // =========================================================================
    assign c[29] = g[28] | (p[28] & c[28]);
    assign c[30] = g[29] | (p[29] & c[29]);
    assign c[31] = g[30] | (p[30] & c[30]);
    assign c[32] = g[31] | (p[31] & c[31]);

    assign block_p[7] = p[28] & p[29] & p[30] & p[31];
    assign block_g[7] = g[31] | (p[31] & g[30]) | (p[31] & p[30] & g[29]) | (p[31] & p[30] & p[29] & g[28]);

    // =========================================================================
    // Second-level carry lookahead (block carries)
    // =========================================================================
    assign block_c[1] = block_g[0] | (block_p[0] & block_c[0]);
    assign block_c[2] = block_g[1] | (block_p[1] & block_c[1]);
    assign block_c[3] = block_g[2] | (block_p[2] & block_c[2]);
    assign block_c[4] = block_g[3] | (block_p[3] & block_c[3]);
    assign block_c[5] = block_g[4] | (block_p[4] & block_c[4]);
    assign block_c[6] = block_g[5] | (block_p[5] & block_c[5]);
    assign block_c[7] = block_g[6] | (block_p[6] & block_c[6]);
    assign block_c[8] = block_g[7] | (block_p[7] & block_c[7]);

    // =========================================================================
    // Final sum generation
    // =========================================================================
    assign sum = p ^ c[31:0];

endmodule